module Total_tcam(input [103:0]key,
input write_clk,
input readen,
input wren,
input resetn,
input [103:0] wr_addr,
input [103:0]rule0,
input [103:0]rule1,
input [103:0]rule2,
input [103:0]rule3,
input [103:0]rule4,
input [103:0]rule5,
input [103:0]rule6,
input [103:0]rule7,
input [103:0]rule8,
input [103:0]rule9,
input [103:0]rule10,
input [103:0]rule11,
input [103:0]rule12,
input [103:0]rule13,
input [103:0]rule14,
input [103:0]rule15,
input [103:0]rule16,
input [103:0]rule17,
input [103:0]rule18,
input [103:0]rule19,
input [103:0]rule20,
input [103:0]rule21,
input [103:0]rule22,
input [103:0]rule23,
input [103:0]rule24,
input [103:0]rule25,
input [103:0]rule26,
input [103:0]rule27,
input [103:0]rule28,
input [103:0]rule29,
input [103:0]rule30,
input [103:0]rule31,
input [103:0]rule32,
input [103:0]rule33,
input [103:0]rule34,
input [103:0]rule35,
input [103:0]rule36,
input [103:0]rule37,
input [103:0]rule38,
input [103:0]rule39,
input [103:0]rule40,
input [103:0]rule41,
input [103:0]rule42,
input [103:0]rule43,
input [103:0]rule44,
input [103:0]rule45,
input [103:0]rule46,
input [103:0]rule47,
input [103:0]rule48,
input [103:0]rule49,
input [103:0]rule50,
input [103:0]rule51,
input [103:0]rule52,
input [103:0]rule53,
input [103:0]rule54,
input [103:0]rule55,
input [103:0]rule56,
input [103:0]rule57,
input [103:0]rule58,
input [103:0]rule59,
input [103:0]rule60,
input [103:0]rule61,
input [103:0]rule62,
input [103:0]rule63,
input [103:0]rule64,
input [103:0]rule65,
input [103:0]rule66,
input [103:0]rule67,
input [103:0]rule68,
input [103:0]rule69,
input [103:0]rule70,
input [103:0]rule71,
input [103:0]rule72,
input [103:0]rule73,
input [103:0]rule74,
input [103:0]rule75,
input [103:0]rule76,
input [103:0]rule77,
input [103:0]rule78,
input [103:0]rule79,
input [103:0]rule80,
input [103:0]rule81,
input [103:0]rule82,
input [103:0]rule83,
input [103:0]rule84,
input [103:0]rule85,
input [103:0]rule86,
input [103:0]rule87,
input [103:0]rule88,
input [103:0]rule89,
input [103:0]rule90,
input [103:0]rule91,
input [103:0]rule92,
input [103:0]rule93,
input [103:0]rule94,
input [103:0]rule95,
input [103:0]rule96,
input [103:0]rule97,
input [103:0]rule98,
input [103:0]rule99,
input [103:0]rule100,
input [103:0]rule101,
input [103:0]rule102,
input [103:0]rule103,
input [103:0]rule104,
input [103:0]rule105,
input [103:0]rule106,
input [103:0]rule107,
input [103:0]rule108,
input [103:0]rule109,
input [103:0]rule110,
input [103:0]rule111,
input [103:0]rule112,
input [103:0]rule113,
input [103:0]rule114,
input [103:0]rule115,
input [103:0]rule116,
input [103:0]rule117,
input [103:0]rule118,
input [103:0]rule119,
output reg [119:0] result);

wire [119:0] data0,data1,data2,data3,data4,data5,data6,data7,data8,data9,data10,data11,data12;
wire [119:0] i_data;
 
Row_of_RAM iRow_of_RAM0(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),
		.rule0(rule0[7:0]),
		.rule1(rule1[7:0]),
		.rule2(rule2[7:0]),
		.rule3(rule3[7:0]),
		.rule4(rule4[7:0]),
		.rule5(rule5[7:0]),
		.rule6(rule6[7:0]),
		.rule7(rule7[7:0]),
		.rule8(rule8[7:0]),
		.rule9(rule9[7:0]),
		.rule10(rule10[7:0]),
		.rule11(rule11[7:0]),
		.rule12(rule12[7:0]),
		.rule13(rule13[7:0]),
		.rule14(rule14[7:0]),
                .rule15(rule15[7:0]),
                .rule16(rule16[7:0]),
                .rule17(rule17[7:0]),
                .rule18(rule18[7:0]),
                .rule19(rule19[7:0]),
                .rule20(rule20[7:0]),
                .rule21(rule21[7:0]),
                .rule22(rule22[7:0]),
                .rule23(rule23[7:0]),
                .rule24(rule24[7:0]),
                .rule25(rule25[7:0]),
                .rule26(rule26[7:0]),
                .rule27(rule27[7:0]),
                .rule28(rule28[7:0]),
                .rule29(rule29[7:0]),
                .rule30(rule30[7:0]),
                .rule31(rule31[7:0]),
                .rule32(rule32[7:0]),
                .rule33(rule33[7:0]),
               	.rule34(rule34[7:0]),
               	.rule35(rule35[7:0]),
                .rule36(rule36[7:0]),
               .rule37(rule37[7:0]),
               .rule38(rule38[7:0]),
               .rule39(rule39[7:0]),
               .rule40(rule40[7:0]),
               .rule41(rule41[7:0]),
               .rule42(rule42[7:0]),
               .rule43(rule43[7:0]),
               .rule44(rule44[7:0]),
               .rule45(rule45[7:0]),
               .rule46(rule46[7:0]),
               .rule47(rule47[7:0]),
               .rule48(rule48[7:0]),
               .rule49(rule49[7:0]),
               .rule50(rule50[7:0]),
               .rule51(rule51[7:0]),
               .rule52(rule52[7:0]),
               .rule53(rule53[7:0]),
               .rule54(rule54[7:0]),
               .rule55(rule55[7:0]),
               .rule56(rule56[7:0]),
               .rule57(rule57[7:0]),
               .rule58(rule58[7:0]),
               .rule59(rule59[7:0]),
               .rule60(rule60[7:0]),
               .rule61(rule61[7:0]),
               .rule62(rule62[7:0]),
               .rule63(rule63[7:0]),
               .rule64(rule64[7:0]),
               .rule65(rule65[7:0]),
               .rule66(rule66[7:0]),
               .rule67(rule67[7:0]),
               .rule68(rule68[7:0]),
               .rule69(rule69[7:0]),
               .rule70(rule70[7:0]),
               .rule71(rule71[7:0]),
               .rule72(rule72[7:0]),
               .rule73(rule73[7:0]),
               .rule74(rule74[7:0]),
               .rule75(rule75[7:0]),
               .rule76(rule76[7:0]),
               .rule77(rule77[7:0]),
               .rule78(rule78[7:0]),
               .rule79(rule79[7:0]),
               .rule80(rule80[7:0]),
               .rule81(rule81[7:0]),
               .rule82(rule82[7:0]),
               .rule83(rule83[7:0]),
               .rule84(rule84[7:0]),
               .rule85(rule85[7:0]),
               .rule86(rule86[7:0]),
               .rule87(rule87[7:0]),
               .rule88(rule88[7:0]),
               .rule89(rule89[7:0]),
               .rule90(rule90[7:0]),
               .rule91(rule91[7:0]),
               .rule92(rule92[7:0]),
               .rule93(rule93[7:0]),
               .rule94(rule94[7:0]),
               .rule95(rule95[7:0]),
               .rule96(rule96[7:0]),
               .rule97(rule97[7:0]),
               .rule98(rule98[7:0]),
               .rule99(rule99[7:0]),
               .rule100(rule100[7:0]),
               .rule101(rule101[7:0]),
               .rule102(rule102[7:0]),
               .rule103(rule103[7:0]),
               .rule104(rule104[7:0]),
               .rule105(rule105[7:0]),
               .rule106(rule106[7:0]),
               .rule107(rule107[7:0]),
               .rule108(rule108[7:0]),
               .rule109(rule109[7:0]),
               .rule110(rule110[7:0]),
               .rule111(rule111[7:0]),
               .rule112(rule112[7:0]),
               .rule113(rule113[7:0]),
               .rule114(rule114[7:0]),
               .rule115(rule115[7:0]),
               .rule116(rule116[7:0]),
               .rule117(rule117[7:0]),
               .rule118(rule118[7:0]),
               .rule119(rule119[7:0]),
		.match(data0));
Row_of_RAM iRow_of_RAM1(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[15:8]),.key(key[15:8]),
		.rule0(rule0[15:8]),
		.rule1(rule1[15:8]),
		.rule2(rule2[15:8]),
		.rule3(rule3[15:8]),
		.rule4(rule4[15:8]),
		.rule5(rule5[15:8]),
		.rule6(rule6[15:8]),
		.rule7(rule7[15:8]),
		.rule8(rule8[15:8]),
		.rule9(rule9[15:8]),
		.rule10(rule10[15:8]),
		.rule11(rule11[15:8]),
		.rule12(rule12[15:8]),
		.rule13(rule13[15:8]),
		.rule14(rule14[15:8]),
                .rule15(rule15[15:8]),
                .rule16(rule16[15:8]),
                .rule17(rule17[15:8]),
                .rule18(rule18[15:8]),
                .rule19(rule19[15:8]),
                .rule20(rule20[15:8]),
                .rule21(rule21[15:8]),
                .rule22(rule22[15:8]),
                .rule23(rule23[15:8]),
                .rule24(rule24[15:8]),
                .rule25(rule25[15:8]),
                .rule26(rule26[15:8]),
                .rule27(rule27[15:8]),
                .rule28(rule28[15:8]),
                .rule29(rule29[15:8]),
                .rule30(rule30[15:8]),
                .rule31(rule31[15:8]),
                .rule32(rule32[15:8]),
                .rule33(rule33[15:8]),
               	.rule34(rule34[15:8]),
               	.rule35(rule35[15:8]),
                .rule36(rule36[15:8]),
               .rule37(rule37[15:8]),
               .rule38(rule38[15:8]),
               .rule39(rule39[15:8]),
               .rule40(rule40[15:8]),
               .rule41(rule41[15:8]),
               .rule42(rule42[15:8]),
               .rule43(rule43[15:8]),
               .rule44(rule44[15:8]),
               .rule45(rule45[15:8]),
               .rule46(rule46[15:8]),
               .rule47(rule47[15:8]),
               .rule48(rule48[15:8]),
               .rule49(rule49[15:8]),
               .rule50(rule50[15:8]),
               .rule51(rule51[15:8]),
               .rule52(rule52[15:8]),
               .rule53(rule53[15:8]),
               .rule54(rule54[15:8]),
               .rule55(rule55[15:8]),
               .rule56(rule56[15:8]),
               .rule57(rule57[15:8]),
               .rule58(rule58[15:8]),
               .rule59(rule59[15:8]),
               .rule60(rule60[15:8]),
               .rule61(rule61[15:8]),
               .rule62(rule62[15:8]),
               .rule63(rule63[15:8]),
               .rule64(rule64[15:8]),
               .rule65(rule65[15:8]),
               .rule66(rule66[15:8]),
               .rule67(rule67[15:8]),
               .rule68(rule68[15:8]),
               .rule69(rule69[15:8]),
               .rule70(rule70[15:8]),
               .rule71(rule71[15:8]),
               .rule72(rule72[15:8]),
               .rule73(rule73[15:8]),
               .rule74(rule74[15:8]),
               .rule75(rule75[15:8]),
               .rule76(rule76[15:8]),
               .rule77(rule77[15:8]),
               .rule78(rule78[15:8]),
               .rule79(rule79[15:8]),
               .rule80(rule80[15:8]),
               .rule81(rule81[15:8]),
               .rule82(rule82[15:8]),
               .rule83(rule83[15:8]),
               .rule84(rule84[15:8]),
               .rule85(rule85[15:8]),
               .rule86(rule86[15:8]),
               .rule87(rule87[15:8]),
               .rule88(rule88[15:8]),
               .rule89(rule89[15:8]),
               .rule90(rule90[15:8]),
               .rule91(rule91[15:8]),
               .rule92(rule92[15:8]),
               .rule93(rule93[15:8]),
               .rule94(rule94[15:8]),
               .rule95(rule95[15:8]),
               .rule96(rule96[15:8]),
               .rule97(rule97[15:8]),
               .rule98(rule98[15:8]),
               .rule99(rule99[15:8]),
               .rule100(rule100[15:8]),
               .rule101(rule101[15:8]),
               .rule102(rule102[15:8]),
               .rule103(rule103[15:8]),
               .rule104(rule104[15:8]),
               .rule105(rule105[15:8]),
               .rule106(rule106[15:8]),
               .rule107(rule107[15:8]),
               .rule108(rule108[15:8]),
               .rule109(rule109[15:8]),
               .rule110(rule110[15:8]),
               .rule111(rule111[15:8]),
               .rule112(rule112[15:8]),
               .rule113(rule113[15:8]),
               .rule114(rule114[15:8]),
               .rule115(rule115[15:8]),
               .rule116(rule116[15:8]),
               .rule117(rule117[15:8]),
               .rule118(rule118[15:8]),
               .rule119(rule119[15:8]),
		.match(data1));
Row_of_RAM iRow_of_RAM2(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[23:16]),.key(key[23:16]),
		.rule0(rule0[23:16]),
		.rule1(rule1[23:16]),
		.rule2(rule2[23:16]),
		.rule3(rule3[23:16]),
		.rule4(rule4[23:16]),
		.rule5(rule5[23:16]),
		.rule6(rule6[23:16]),
		.rule7(rule7[23:16]),
		.rule8(rule8[23:16]),
		.rule9(rule9[23:16]),
		.rule10(rule10[23:16]),
		.rule11(rule11[23:16]),
		.rule12(rule12[23:16]),
		.rule13(rule13[23:16]),
		.rule14(rule14[23:16]),
                .rule15(rule15[23:16]),
                .rule16(rule16[23:16]),
                .rule17(rule17[23:16]),
                .rule18(rule18[23:16]),
                .rule19(rule19[23:16]),
                .rule20(rule20[23:16]),
                .rule21(rule21[23:16]),
                .rule22(rule22[23:16]),
                .rule23(rule23[23:16]),
                .rule24(rule24[23:16]),
                .rule25(rule25[23:16]),
                .rule26(rule26[23:16]),
                .rule27(rule27[23:16]),
                .rule28(rule28[23:16]),
                .rule29(rule29[23:16]),
                .rule30(rule30[23:16]),
                .rule31(rule31[23:16]),
                .rule32(rule32[23:16]),
                .rule33(rule33[23:16]),
               	.rule34(rule34[23:16]),
               	.rule35(rule35[23:16]),
                .rule36(rule36[23:16]),
               .rule37(rule37[23:16]),
               .rule38(rule38[23:16]),
               .rule39(rule39[23:16]),
               .rule40(rule40[23:16]),
               .rule41(rule41[23:16]),
               .rule42(rule42[23:16]),
               .rule43(rule43[23:16]),
               .rule44(rule44[23:16]),
               .rule45(rule45[23:16]),
               .rule46(rule46[23:16]),
               .rule47(rule47[23:16]),
               .rule48(rule48[23:16]),
               .rule49(rule49[23:16]),
               .rule50(rule50[23:16]),
               .rule51(rule51[23:16]),
               .rule52(rule52[23:16]),
               .rule53(rule53[23:16]),
               .rule54(rule54[23:16]),
               .rule55(rule55[23:16]),
               .rule56(rule56[23:16]),
               .rule57(rule57[23:16]),
               .rule58(rule58[23:16]),
               .rule59(rule59[23:16]),
               .rule60(rule60[23:16]),
               .rule61(rule61[23:16]),
               .rule62(rule62[23:16]),
               .rule63(rule63[23:16]),
               .rule64(rule64[23:16]),
               .rule65(rule65[23:16]),
               .rule66(rule66[23:16]),
               .rule67(rule67[23:16]),
               .rule68(rule68[23:16]),
               .rule69(rule69[23:16]),
               .rule70(rule70[23:16]),
               .rule71(rule71[23:16]),
               .rule72(rule72[23:16]),
               .rule73(rule73[23:16]),
               .rule74(rule74[23:16]),
               .rule75(rule75[23:16]),
               .rule76(rule76[23:16]),
               .rule77(rule77[23:16]),
               .rule78(rule78[23:16]),
               .rule79(rule79[23:16]),
               .rule80(rule80[23:16]),
               .rule81(rule81[23:16]),
               .rule82(rule82[23:16]),
               .rule83(rule83[23:16]),
               .rule84(rule84[23:16]),
               .rule85(rule85[23:16]),
               .rule86(rule86[23:16]),
               .rule87(rule87[23:16]),
               .rule88(rule88[23:16]),
               .rule89(rule89[23:16]),
               .rule90(rule90[23:16]),
               .rule91(rule91[23:16]),
               .rule92(rule92[23:16]),
               .rule93(rule93[23:16]),
               .rule94(rule94[23:16]),
               .rule95(rule95[23:16]),
               .rule96(rule96[23:16]),
               .rule97(rule97[23:16]),
               .rule98(rule98[23:16]),
               .rule99(rule99[23:16]),
               .rule100(rule100[23:16]),
               .rule101(rule101[23:16]),
               .rule102(rule102[23:16]),
               .rule103(rule103[23:16]),
               .rule104(rule104[23:16]),
               .rule105(rule105[23:16]),
               .rule106(rule106[23:16]),
               .rule107(rule107[23:16]),
               .rule108(rule108[23:16]),
               .rule109(rule109[23:16]),
               .rule110(rule110[23:16]),
               .rule111(rule111[23:16]),
               .rule112(rule112[23:16]),
               .rule113(rule113[23:16]),
               .rule114(rule114[23:16]),
               .rule115(rule115[23:16]),
               .rule116(rule116[23:16]),
               .rule117(rule117[23:16]),
               .rule118(rule118[23:16]),
               .rule119(rule119[23:16]),
		.match(data2));
Row_of_RAM iRow_of_RAM3(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[31:24]),.key(key[31:24]),
		.rule0(rule0[31:24]),
		.rule1(rule1[31:24]),
		.rule2(rule2[31:24]),
		.rule3(rule3[31:24]),
		.rule4(rule4[31:24]),
		.rule5(rule5[31:24]),
		.rule6(rule6[31:24]),
		.rule7(rule7[31:24]),
		.rule8(rule8[31:24]),
		.rule9(rule9[31:24]),
		.rule10(rule10[31:24]),
		.rule11(rule11[31:24]),
		.rule12(rule12[31:24]),
		.rule13(rule13[31:24]),
		.rule14(rule14[31:24]),
                .rule15(rule15[31:24]),
                .rule16(rule16[31:24]),
                .rule17(rule17[31:24]),
                .rule18(rule18[31:24]),
                .rule19(rule19[31:24]),
                .rule20(rule20[31:24]),
                .rule21(rule21[31:24]),
                .rule22(rule22[31:24]),
                .rule23(rule23[31:24]),
                .rule24(rule24[31:24]),
                .rule25(rule25[31:24]),
                .rule26(rule26[31:24]),
                .rule27(rule27[31:24]),
                .rule28(rule28[31:24]),
                .rule29(rule29[31:24]),
                .rule30(rule30[31:24]),
                .rule31(rule31[31:24]),
                .rule32(rule32[31:24]),
                .rule33(rule33[31:24]),
               	.rule34(rule34[31:24]),
               	.rule35(rule35[31:24]),
                .rule36(rule36[31:24]),
               .rule37(rule37[31:24]),
               .rule38(rule38[31:24]),
               .rule39(rule39[31:24]),
               .rule40(rule40[31:24]),
               .rule41(rule41[31:24]),
               .rule42(rule42[31:24]),
               .rule43(rule43[31:24]),
               .rule44(rule44[31:24]),
               .rule45(rule45[31:24]),
               .rule46(rule46[31:24]),
               .rule47(rule47[31:24]),
               .rule48(rule48[31:24]),
               .rule49(rule49[31:24]),
               .rule50(rule50[31:24]),
               .rule51(rule51[31:24]),
               .rule52(rule52[31:24]),
               .rule53(rule53[31:24]),
               .rule54(rule54[31:24]),
               .rule55(rule55[31:24]),
               .rule56(rule56[31:24]),
               .rule57(rule57[31:24]),
               .rule58(rule58[31:24]),
               .rule59(rule59[31:24]),
               .rule60(rule60[31:24]),
               .rule61(rule61[31:24]),
               .rule62(rule62[31:24]),
               .rule63(rule63[31:24]),
               .rule64(rule64[31:24]),
               .rule65(rule65[31:24]),
               .rule66(rule66[31:24]),
               .rule67(rule67[31:24]),
               .rule68(rule68[31:24]),
               .rule69(rule69[31:24]),
               .rule70(rule70[31:24]),
               .rule71(rule71[31:24]),
               .rule72(rule72[31:24]),
               .rule73(rule73[31:24]),
               .rule74(rule74[31:24]),
               .rule75(rule75[31:24]),
               .rule76(rule76[31:24]),
               .rule77(rule77[31:24]),
               .rule78(rule78[31:24]),
               .rule79(rule79[31:24]),
               .rule80(rule80[31:24]),
               .rule81(rule81[31:24]),
               .rule82(rule82[31:24]),
               .rule83(rule83[31:24]),
               .rule84(rule84[31:24]),
               .rule85(rule85[31:24]),
               .rule86(rule86[31:24]),
               .rule87(rule87[31:24]),
               .rule88(rule88[31:24]),
               .rule89(rule89[31:24]),
               .rule90(rule90[31:24]),
               .rule91(rule91[31:24]),
               .rule92(rule92[31:24]),
               .rule93(rule93[31:24]),
               .rule94(rule94[31:24]),
               .rule95(rule95[31:24]),
               .rule96(rule96[31:24]),
               .rule97(rule97[31:24]),
               .rule98(rule98[31:24]),
               .rule99(rule99[31:24]),
               .rule100(rule100[31:24]),
               .rule101(rule101[31:24]),
               .rule102(rule102[31:24]),
               .rule103(rule103[31:24]),
               .rule104(rule104[31:24]),
               .rule105(rule105[31:24]),
               .rule106(rule106[31:24]),
               .rule107(rule107[31:24]),
               .rule108(rule108[31:24]),
               .rule109(rule109[31:24]),
               .rule110(rule110[31:24]),
               .rule111(rule111[31:24]),
               .rule112(rule112[31:24]),
               .rule113(rule113[31:24]),
               .rule114(rule114[31:24]),
               .rule115(rule115[31:24]),
               .rule116(rule116[31:24]),
               .rule117(rule117[31:24]),
               .rule118(rule118[31:24]),
               .rule119(rule119[31:24]),
		.match(data3));
Row_of_RAM iRow_of_RAM4(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[39:32]),.key(key[39:32]),
		.rule0(rule0[39:32]),
		.rule1(rule1[39:32]),
		.rule2(rule2[39:32]),
		.rule3(rule3[39:32]),
		.rule4(rule4[39:32]),
		.rule5(rule5[39:32]),
		.rule6(rule6[39:32]),
		.rule7(rule7[39:32]),
		.rule8(rule8[39:32]),
		.rule9(rule9[39:32]),
		.rule10(rule10[39:32]),
		.rule11(rule11[39:32]),
		.rule12(rule12[39:32]),
		.rule13(rule13[39:32]),
		.rule14(rule14[39:32]),
                .rule15(rule15[39:32]),
                .rule16(rule16[39:32]),
                .rule17(rule17[39:32]),
                .rule18(rule18[39:32]),
                .rule19(rule19[39:32]),
                .rule20(rule20[39:32]),
                .rule21(rule21[39:32]),
                .rule22(rule22[39:32]),
                .rule23(rule23[39:32]),
                .rule24(rule24[39:32]),
                .rule25(rule25[39:32]),
                .rule26(rule26[39:32]),
                .rule27(rule27[39:32]),
                .rule28(rule28[39:32]),
                .rule29(rule29[39:32]),
                .rule30(rule30[39:32]),
                .rule31(rule31[39:32]),
                .rule32(rule32[39:32]),
                .rule33(rule33[39:32]),
               	.rule34(rule34[39:32]),
               	.rule35(rule35[39:32]),
                .rule36(rule36[39:32]),
               .rule37(rule37[39:32]),
               .rule38(rule38[39:32]),
               .rule39(rule39[39:32]),
               .rule40(rule40[39:32]),
               .rule41(rule41[39:32]),
               .rule42(rule42[39:32]),
               .rule43(rule43[39:32]),
               .rule44(rule44[39:32]),
               .rule45(rule45[39:32]),
               .rule46(rule46[39:32]),
               .rule47(rule47[39:32]),
               .rule48(rule48[39:32]),
               .rule49(rule49[39:32]),
               .rule50(rule50[39:32]),
               .rule51(rule51[39:32]),
               .rule52(rule52[39:32]),
               .rule53(rule53[39:32]),
               .rule54(rule54[39:32]),
               .rule55(rule55[39:32]),
               .rule56(rule56[39:32]),
               .rule57(rule57[39:32]),
               .rule58(rule58[39:32]),
               .rule59(rule59[39:32]),
               .rule60(rule60[39:32]),
               .rule61(rule61[39:32]),
               .rule62(rule62[39:32]),
               .rule63(rule63[39:32]),
               .rule64(rule64[39:32]),
               .rule65(rule65[39:32]),
               .rule66(rule66[39:32]),
               .rule67(rule67[39:32]),
               .rule68(rule68[39:32]),
               .rule69(rule69[39:32]),
               .rule70(rule70[39:32]),
               .rule71(rule71[39:32]),
               .rule72(rule72[39:32]),
               .rule73(rule73[39:32]),
               .rule74(rule74[39:32]),
               .rule75(rule75[39:32]),
               .rule76(rule76[39:32]),
               .rule77(rule77[39:32]),
               .rule78(rule78[39:32]),
               .rule79(rule79[39:32]),
               .rule80(rule80[39:32]),
               .rule81(rule81[39:32]),
               .rule82(rule82[39:32]),
               .rule83(rule83[39:32]),
               .rule84(rule84[39:32]),
               .rule85(rule85[39:32]),
               .rule86(rule86[39:32]),
               .rule87(rule87[39:32]),
               .rule88(rule88[39:32]),
               .rule89(rule89[39:32]),
               .rule90(rule90[39:32]),
               .rule91(rule91[39:32]),
               .rule92(rule92[39:32]),
               .rule93(rule93[39:32]),
               .rule94(rule94[39:32]),
               .rule95(rule95[39:32]),
               .rule96(rule96[39:32]),
               .rule97(rule97[39:32]),
               .rule98(rule98[39:32]),
               .rule99(rule99[39:32]),
               .rule100(rule100[39:32]),
               .rule101(rule101[39:32]),
               .rule102(rule102[39:32]),
               .rule103(rule103[39:32]),
               .rule104(rule104[39:32]),
               .rule105(rule105[39:32]),
               .rule106(rule106[39:32]),
               .rule107(rule107[39:32]),
               .rule108(rule108[39:32]),
               .rule109(rule109[39:32]),
               .rule110(rule110[39:32]),
               .rule111(rule111[39:32]),
               .rule112(rule112[39:32]),
               .rule113(rule113[39:32]),
               .rule114(rule114[39:32]),
               .rule115(rule115[39:32]),
               .rule116(rule116[39:32]),
               .rule117(rule117[39:32]),
               .rule118(rule118[39:32]),
               .rule119(rule119[39:32]),
		.match(data4));
Row_of_RAM iRow_of_RAM5(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[47:40]),.key(key[47:40]),
		.rule0(rule0[47:40]),
		.rule1(rule1[47:40]),
		.rule2(rule2[47:40]),
		.rule3(rule3[47:40]),
		.rule4(rule4[47:40]),
		.rule5(rule5[47:40]),
		.rule6(rule6[47:40]),
		.rule7(rule7[47:40]),
		.rule8(rule8[47:40]),
		.rule9(rule9[47:40]),
		.rule10(rule10[47:40]),
		.rule11(rule11[47:40]),
		.rule12(rule12[47:40]),
		.rule13(rule13[47:40]),
		.rule14(rule14[47:40]),
                .rule15(rule15[47:40]),
                .rule16(rule16[47:40]),
                .rule17(rule17[47:40]),
                .rule18(rule18[47:40]),
                .rule19(rule19[47:40]),
                .rule20(rule20[47:40]),
                .rule21(rule21[47:40]),
                .rule22(rule22[47:40]),
                .rule23(rule23[47:40]),
                .rule24(rule24[47:40]),
                .rule25(rule25[47:40]),
                .rule26(rule26[47:40]),
                .rule27(rule27[47:40]),
                .rule28(rule28[47:40]),
                .rule29(rule29[47:40]),
                .rule30(rule30[47:40]),
                .rule31(rule31[47:40]),
                .rule32(rule32[47:40]),
                .rule33(rule33[47:40]),
               	.rule34(rule34[47:40]),
               	.rule35(rule35[47:40]),
                .rule36(rule36[47:40]),
               .rule37(rule37[47:40]),
               .rule38(rule38[47:40]),
               .rule39(rule39[47:40]),
               .rule40(rule40[47:40]),
               .rule41(rule41[47:40]),
               .rule42(rule42[47:40]),
               .rule43(rule43[47:40]),
               .rule44(rule44[47:40]),
               .rule45(rule45[47:40]),
               .rule46(rule46[47:40]),
               .rule47(rule47[47:40]),
               .rule48(rule48[47:40]),
               .rule49(rule49[47:40]),
               .rule50(rule50[47:40]),
               .rule51(rule51[47:40]),
               .rule52(rule52[47:40]),
               .rule53(rule53[47:40]),
               .rule54(rule54[47:40]),
               .rule55(rule55[47:40]),
               .rule56(rule56[47:40]),
               .rule57(rule57[47:40]),
               .rule58(rule58[47:40]),
               .rule59(rule59[47:40]),
               .rule60(rule60[47:40]),
               .rule61(rule61[47:40]),
               .rule62(rule62[47:40]),
               .rule63(rule63[47:40]),
               .rule64(rule64[47:40]),
               .rule65(rule65[47:40]),
               .rule66(rule66[47:40]),
               .rule67(rule67[47:40]),
               .rule68(rule68[47:40]),
               .rule69(rule69[47:40]),
               .rule70(rule70[47:40]),
               .rule71(rule71[47:40]),
               .rule72(rule72[47:40]),
               .rule73(rule73[47:40]),
               .rule74(rule74[47:40]),
               .rule75(rule75[47:40]),
               .rule76(rule76[47:40]),
               .rule77(rule77[47:40]),
               .rule78(rule78[47:40]),
               .rule79(rule79[47:40]),
               .rule80(rule80[47:40]),
               .rule81(rule81[47:40]),
               .rule82(rule82[47:40]),
               .rule83(rule83[47:40]),
               .rule84(rule84[47:40]),
               .rule85(rule85[47:40]),
               .rule86(rule86[47:40]),
               .rule87(rule87[47:40]),
               .rule88(rule88[47:40]),
               .rule89(rule89[47:40]),
               .rule90(rule90[47:40]),
               .rule91(rule91[47:40]),
               .rule92(rule92[47:40]),
               .rule93(rule93[47:40]),
               .rule94(rule94[47:40]),
               .rule95(rule95[47:40]),
               .rule96(rule96[47:40]),
               .rule97(rule97[47:40]),
               .rule98(rule98[47:40]),
               .rule99(rule99[47:40]),
               .rule100(rule100[47:40]),
               .rule101(rule101[47:40]),
               .rule102(rule102[47:40]),
               .rule103(rule103[47:40]),
               .rule104(rule104[47:40]),
               .rule105(rule105[47:40]),
               .rule106(rule106[47:40]),
               .rule107(rule107[47:40]),
               .rule108(rule108[47:40]),
               .rule109(rule109[47:40]),
               .rule110(rule110[47:40]),
               .rule111(rule111[47:40]),
               .rule112(rule112[47:40]),
               .rule113(rule113[47:40]),
               .rule114(rule114[47:40]),
               .rule115(rule115[47:40]),
               .rule116(rule116[47:40]),
               .rule117(rule117[47:40]),
               .rule118(rule118[47:40]),
               .rule119(rule119[47:40]),
		.match(data5));
Row_of_RAM iRow_of_RAM6(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[55:48]),.key(key[55:48]),
		.rule0(rule0[55:48]),
		.rule1(rule1[55:48]),
		.rule2(rule2[55:48]),
		.rule3(rule3[55:48]),
		.rule4(rule4[55:48]),
		.rule5(rule5[55:48]),
		.rule6(rule6[55:48]),
		.rule7(rule7[55:48]),
		.rule8(rule8[55:48]),
		.rule9(rule9[55:48]),
		.rule10(rule10[55:48]),
		.rule11(rule11[55:48]),
		.rule12(rule12[55:48]),
		.rule13(rule13[55:48]),
		.rule14(rule14[55:48]),
                .rule15(rule15[55:48]),
                .rule16(rule16[55:48]),
                .rule17(rule17[55:48]),
                .rule18(rule18[55:48]),
                .rule19(rule19[55:48]),
                .rule20(rule20[55:48]),
                .rule21(rule21[55:48]),
                .rule22(rule22[55:48]),
                .rule23(rule23[55:48]),
                .rule24(rule24[55:48]),
                .rule25(rule25[55:48]),
                .rule26(rule26[55:48]),
                .rule27(rule27[55:48]),
                .rule28(rule28[55:48]),
                .rule29(rule29[55:48]),
                .rule30(rule30[55:48]),
                .rule31(rule31[55:48]),
                .rule32(rule32[55:48]),
                .rule33(rule33[55:48]),
               	.rule34(rule34[55:48]),
               	.rule35(rule35[55:48]),
                .rule36(rule36[55:48]),
               .rule37(rule37[55:48]),
               .rule38(rule38[55:48]),
               .rule39(rule39[55:48]),
               .rule40(rule40[55:48]),
               .rule41(rule41[55:48]),
               .rule42(rule42[55:48]),
               .rule43(rule43[55:48]),
               .rule44(rule44[55:48]),
               .rule45(rule45[55:48]),
               .rule46(rule46[55:48]),
               .rule47(rule47[55:48]),
               .rule48(rule48[55:48]),
               .rule49(rule49[55:48]),
               .rule50(rule50[55:48]),
               .rule51(rule51[55:48]),
               .rule52(rule52[55:48]),
               .rule53(rule53[55:48]),
               .rule54(rule54[55:48]),
               .rule55(rule55[55:48]),
               .rule56(rule56[55:48]),
               .rule57(rule57[55:48]),
               .rule58(rule58[55:48]),
               .rule59(rule59[55:48]),
               .rule60(rule60[55:48]),
               .rule61(rule61[55:48]),
               .rule62(rule62[55:48]),
               .rule63(rule63[55:48]),
               .rule64(rule64[55:48]),
               .rule65(rule65[55:48]),
               .rule66(rule66[55:48]),
               .rule67(rule67[55:48]),
               .rule68(rule68[55:48]),
               .rule69(rule69[55:48]),
               .rule70(rule70[55:48]),
               .rule71(rule71[55:48]),
               .rule72(rule72[55:48]),
               .rule73(rule73[55:48]),
               .rule74(rule74[55:48]),
               .rule75(rule75[55:48]),
               .rule76(rule76[55:48]),
               .rule77(rule77[55:48]),
               .rule78(rule78[55:48]),
               .rule79(rule79[55:48]),
               .rule80(rule80[55:48]),
               .rule81(rule81[55:48]),
               .rule82(rule82[55:48]),
               .rule83(rule83[55:48]),
               .rule84(rule84[55:48]),
               .rule85(rule85[55:48]),
               .rule86(rule86[55:48]),
               .rule87(rule87[55:48]),
               .rule88(rule88[55:48]),
               .rule89(rule89[55:48]),
               .rule90(rule90[55:48]),
               .rule91(rule91[55:48]),
               .rule92(rule92[55:48]),
               .rule93(rule93[55:48]),
               .rule94(rule94[55:48]),
               .rule95(rule95[55:48]),
               .rule96(rule96[55:48]),
               .rule97(rule97[55:48]),
               .rule98(rule98[55:48]),
               .rule99(rule99[55:48]),
               .rule100(rule100[55:48]),
               .rule101(rule101[55:48]),
               .rule102(rule102[55:48]),
               .rule103(rule103[55:48]),
               .rule104(rule104[55:48]),
               .rule105(rule105[55:48]),
               .rule106(rule106[55:48]),
               .rule107(rule107[55:48]),
               .rule108(rule108[55:48]),
               .rule109(rule109[55:48]),
               .rule110(rule110[55:48]),
               .rule111(rule111[55:48]),
               .rule112(rule112[55:48]),
               .rule113(rule113[55:48]),
               .rule114(rule114[55:48]),
               .rule115(rule115[55:48]),
               .rule116(rule116[55:48]),
               .rule117(rule117[55:48]),
               .rule118(rule118[55:48]),
               .rule119(rule119[55:48]),
		.match(data6));
Row_of_RAM iRow_of_RAM7(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[63:56]),.key(key[63:56]),
		.rule0(rule0[63:56]),
		.rule1(rule1[63:56]),
		.rule2(rule2[63:56]),
		.rule3(rule3[63:56]),
		.rule4(rule4[63:56]),
		.rule5(rule5[63:56]),
		.rule6(rule6[63:56]),
		.rule7(rule7[63:56]),
		.rule8(rule8[63:56]),
		.rule9(rule9[63:56]),
		.rule10(rule10[63:56]),
		.rule11(rule11[63:56]),
		.rule12(rule12[63:56]),
		.rule13(rule13[63:56]),
		.rule14(rule14[63:56]),
                .rule15(rule15[63:56]),
                .rule16(rule16[63:56]),
                .rule17(rule17[63:56]),
                .rule18(rule18[63:56]),
                .rule19(rule19[63:56]),
                .rule20(rule20[63:56]),
                .rule21(rule21[63:56]),
                .rule22(rule22[63:56]),
                .rule23(rule23[63:56]),
                .rule24(rule24[63:56]),
                .rule25(rule25[63:56]),
                .rule26(rule26[63:56]),
                .rule27(rule27[63:56]),
                .rule28(rule28[63:56]),
                .rule29(rule29[63:56]),
                .rule30(rule30[63:56]),
                .rule31(rule31[63:56]),
                .rule32(rule32[63:56]),
                .rule33(rule33[63:56]),
               	.rule34(rule34[63:56]),
               	.rule35(rule35[63:56]),
                .rule36(rule36[63:56]),
               .rule37(rule37[63:56]),
               .rule38(rule38[63:56]),
               .rule39(rule39[63:56]),
               .rule40(rule40[63:56]),
               .rule41(rule41[63:56]),
               .rule42(rule42[63:56]),
               .rule43(rule43[63:56]),
               .rule44(rule44[63:56]),
               .rule45(rule45[63:56]),
               .rule46(rule46[63:56]),
               .rule47(rule47[63:56]),
               .rule48(rule48[63:56]),
               .rule49(rule49[63:56]),
               .rule50(rule50[63:56]),
               .rule51(rule51[63:56]),
               .rule52(rule52[63:56]),
               .rule53(rule53[63:56]),
               .rule54(rule54[63:56]),
               .rule55(rule55[63:56]),
               .rule56(rule56[63:56]),
               .rule57(rule57[63:56]),
               .rule58(rule58[63:56]),
               .rule59(rule59[63:56]),
               .rule60(rule60[63:56]),
               .rule61(rule61[63:56]),
               .rule62(rule62[63:56]),
               .rule63(rule63[63:56]),
               .rule64(rule64[63:56]),
               .rule65(rule65[63:56]),
               .rule66(rule66[63:56]),
               .rule67(rule67[63:56]),
               .rule68(rule68[63:56]),
               .rule69(rule69[63:56]),
               .rule70(rule70[63:56]),
               .rule71(rule71[63:56]),
               .rule72(rule72[63:56]),
               .rule73(rule73[63:56]),
               .rule74(rule74[63:56]),
               .rule75(rule75[63:56]),
               .rule76(rule76[63:56]),
               .rule77(rule77[63:56]),
               .rule78(rule78[63:56]),
               .rule79(rule79[63:56]),
               .rule80(rule80[63:56]),
               .rule81(rule81[63:56]),
               .rule82(rule82[63:56]),
               .rule83(rule83[63:56]),
               .rule84(rule84[63:56]),
               .rule85(rule85[63:56]),
               .rule86(rule86[63:56]),
               .rule87(rule87[63:56]),
               .rule88(rule88[63:56]),
               .rule89(rule89[63:56]),
               .rule90(rule90[63:56]),
               .rule91(rule91[63:56]),
               .rule92(rule92[63:56]),
               .rule93(rule93[63:56]),
               .rule94(rule94[63:56]),
               .rule95(rule95[63:56]),
               .rule96(rule96[63:56]),
               .rule97(rule97[63:56]),
               .rule98(rule98[63:56]),
               .rule99(rule99[63:56]),
               .rule100(rule100[63:56]),
               .rule101(rule101[63:56]),
               .rule102(rule102[63:56]),
               .rule103(rule103[63:56]),
               .rule104(rule104[63:56]),
               .rule105(rule105[63:56]),
               .rule106(rule106[63:56]),
               .rule107(rule107[63:56]),
               .rule108(rule108[63:56]),
               .rule109(rule109[63:56]),
               .rule110(rule110[63:56]),
               .rule111(rule111[63:56]),
               .rule112(rule112[63:56]),
               .rule113(rule113[63:56]),
               .rule114(rule114[63:56]),
               .rule115(rule115[63:56]),
               .rule116(rule116[63:56]),
               .rule117(rule117[63:56]),
               .rule118(rule118[63:56]),
               .rule119(rule119[63:56]),
		.match(data7));
Row_of_RAM iRow_of_RAM8(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[71:64]),.key(key[71:64]),
		.rule0(rule0[71:64]),
		.rule1(rule1[71:64]),
		.rule2(rule2[71:64]),
		.rule3(rule3[71:64]),
		.rule4(rule4[71:64]),
		.rule5(rule5[71:64]),
		.rule6(rule6[71:64]),
		.rule7(rule7[71:64]),
		.rule8(rule8[71:64]),
		.rule9(rule9[71:64]),
		.rule10(rule10[71:64]),
		.rule11(rule11[71:64]),
		.rule12(rule12[71:64]),
		.rule13(rule13[71:64]),
		.rule14(rule14[71:64]),
                .rule15(rule15[71:64]),
                .rule16(rule16[71:64]),
                .rule17(rule17[71:64]),
                .rule18(rule18[71:64]),
                .rule19(rule19[71:64]),
                .rule20(rule20[71:64]),
                .rule21(rule21[71:64]),
                .rule22(rule22[71:64]),
                .rule23(rule23[71:64]),
                .rule24(rule24[71:64]),
                .rule25(rule25[71:64]),
                .rule26(rule26[71:64]),
                .rule27(rule27[71:64]),
                .rule28(rule28[71:64]),
                .rule29(rule29[71:64]),
                .rule30(rule30[71:64]),
                .rule31(rule31[71:64]),
                .rule32(rule32[71:64]),
                .rule33(rule33[71:64]),
               	.rule34(rule34[71:64]),
               	.rule35(rule35[71:64]),
                .rule36(rule36[71:64]),
               .rule37(rule37[71:64]),
               .rule38(rule38[71:64]),
               .rule39(rule39[71:64]),
               .rule40(rule40[71:64]),
               .rule41(rule41[71:64]),
               .rule42(rule42[71:64]),
               .rule43(rule43[71:64]),
               .rule44(rule44[71:64]),
               .rule45(rule45[71:64]),
               .rule46(rule46[71:64]),
               .rule47(rule47[71:64]),
               .rule48(rule48[71:64]),
               .rule49(rule49[71:64]),
               .rule50(rule50[71:64]),
               .rule51(rule51[71:64]),
               .rule52(rule52[71:64]),
               .rule53(rule53[71:64]),
               .rule54(rule54[71:64]),
               .rule55(rule55[71:64]),
               .rule56(rule56[71:64]),
               .rule57(rule57[71:64]),
               .rule58(rule58[71:64]),
               .rule59(rule59[71:64]),
               .rule60(rule60[71:64]),
               .rule61(rule61[71:64]),
               .rule62(rule62[71:64]),
               .rule63(rule63[71:64]),
               .rule64(rule64[71:64]),
               .rule65(rule65[71:64]),
               .rule66(rule66[71:64]),
               .rule67(rule67[71:64]),
               .rule68(rule68[71:64]),
               .rule69(rule69[71:64]),
               .rule70(rule70[71:64]),
               .rule71(rule71[71:64]),
               .rule72(rule72[71:64]),
               .rule73(rule73[71:64]),
               .rule74(rule74[71:64]),
               .rule75(rule75[71:64]),
               .rule76(rule76[71:64]),
               .rule77(rule77[71:64]),
               .rule78(rule78[71:64]),
               .rule79(rule79[71:64]),
               .rule80(rule80[71:64]),
               .rule81(rule81[71:64]),
               .rule82(rule82[71:64]),
               .rule83(rule83[71:64]),
               .rule84(rule84[71:64]),
               .rule85(rule85[71:64]),
               .rule86(rule86[71:64]),
               .rule87(rule87[71:64]),
               .rule88(rule88[71:64]),
               .rule89(rule89[71:64]),
               .rule90(rule90[71:64]),
               .rule91(rule91[71:64]),
               .rule92(rule92[71:64]),
               .rule93(rule93[71:64]),
               .rule94(rule94[71:64]),
               .rule95(rule95[71:64]),
               .rule96(rule96[71:64]),
               .rule97(rule97[71:64]),
               .rule98(rule98[71:64]),
               .rule99(rule99[71:64]),
               .rule100(rule100[71:64]),
               .rule101(rule101[71:64]),
               .rule102(rule102[71:64]),
               .rule103(rule103[71:64]),
               .rule104(rule104[71:64]),
               .rule105(rule105[71:64]),
               .rule106(rule106[71:64]),
               .rule107(rule107[71:64]),
               .rule108(rule108[71:64]),
               .rule109(rule109[71:64]),
               .rule110(rule110[71:64]),
               .rule111(rule111[71:64]),
               .rule112(rule112[71:64]),
               .rule113(rule113[71:64]),
               .rule114(rule114[71:64]),
               .rule115(rule115[71:64]),
               .rule116(rule116[71:64]),
               .rule117(rule117[71:64]),
               .rule118(rule118[71:64]),
               .rule119(rule119[71:64]),
		.match(data8));
Row_of_RAM iRow_of_RAM9(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[79:72]),.key(key[79:72]),
		.rule0(rule0[79:72]),
		.rule1(rule1[79:72]),
		.rule2(rule2[79:72]),
		.rule3(rule3[79:72]),
		.rule4(rule4[79:72]),
		.rule5(rule5[79:72]),
		.rule6(rule6[79:72]),
		.rule7(rule7[79:72]),
		.rule8(rule8[79:72]),
		.rule9(rule9[79:72]),
		.rule10(rule10[79:72]),
		.rule11(rule11[79:72]),
		.rule12(rule12[79:72]),
		.rule13(rule13[79:72]),
		.rule14(rule14[79:72]),
                .rule15(rule15[79:72]),
                .rule16(rule16[79:72]),
                .rule17(rule17[79:72]),
                .rule18(rule18[79:72]),
                .rule19(rule19[79:72]),
                .rule20(rule20[79:72]),
                .rule21(rule21[79:72]),
                .rule22(rule22[79:72]),
                .rule23(rule23[79:72]),
                .rule24(rule24[79:72]),
                .rule25(rule25[79:72]),
                .rule26(rule26[79:72]),
                .rule27(rule27[79:72]),
                .rule28(rule28[79:72]),
                .rule29(rule29[79:72]),
                .rule30(rule30[79:72]),
                .rule31(rule31[79:72]),
                .rule32(rule32[79:72]),
                .rule33(rule33[79:72]),
               	.rule34(rule34[79:72]),
               	.rule35(rule35[79:72]),
                .rule36(rule36[79:72]),
               .rule37(rule37[79:72]),
               .rule38(rule38[79:72]),
               .rule39(rule39[79:72]),
               .rule40(rule40[79:72]),
               .rule41(rule41[79:72]),
               .rule42(rule42[79:72]),
               .rule43(rule43[79:72]),
               .rule44(rule44[79:72]),
               .rule45(rule45[79:72]),
               .rule46(rule46[79:72]),
               .rule47(rule47[79:72]),
               .rule48(rule48[79:72]),
               .rule49(rule49[79:72]),
               .rule50(rule50[79:72]),
               .rule51(rule51[79:72]),
               .rule52(rule52[79:72]),
               .rule53(rule53[79:72]),
               .rule54(rule54[79:72]),
               .rule55(rule55[79:72]),
               .rule56(rule56[79:72]),
               .rule57(rule57[79:72]),
               .rule58(rule58[79:72]),
               .rule59(rule59[79:72]),
               .rule60(rule60[79:72]),
               .rule61(rule61[79:72]),
               .rule62(rule62[79:72]),
               .rule63(rule63[79:72]),
               .rule64(rule64[79:72]),
               .rule65(rule65[79:72]),
               .rule66(rule66[79:72]),
               .rule67(rule67[79:72]),
               .rule68(rule68[79:72]),
               .rule69(rule69[79:72]),
               .rule70(rule70[79:72]),
               .rule71(rule71[79:72]),
               .rule72(rule72[79:72]),
               .rule73(rule73[79:72]),
               .rule74(rule74[79:72]),
               .rule75(rule75[79:72]),
               .rule76(rule76[79:72]),
               .rule77(rule77[79:72]),
               .rule78(rule78[79:72]),
               .rule79(rule79[79:72]),
               .rule80(rule80[79:72]),
               .rule81(rule81[79:72]),
               .rule82(rule82[79:72]),
               .rule83(rule83[79:72]),
               .rule84(rule84[79:72]),
               .rule85(rule85[79:72]),
               .rule86(rule86[79:72]),
               .rule87(rule87[79:72]),
               .rule88(rule88[79:72]),
               .rule89(rule89[79:72]),
               .rule90(rule90[79:72]),
               .rule91(rule91[79:72]),
               .rule92(rule92[79:72]),
               .rule93(rule93[79:72]),
               .rule94(rule94[79:72]),
               .rule95(rule95[79:72]),
               .rule96(rule96[79:72]),
               .rule97(rule97[79:72]),
               .rule98(rule98[79:72]),
               .rule99(rule99[79:72]),
               .rule100(rule100[79:72]),
               .rule101(rule101[79:72]),
               .rule102(rule102[79:72]),
               .rule103(rule103[79:72]),
               .rule104(rule104[79:72]),
               .rule105(rule105[79:72]),
               .rule106(rule106[79:72]),
               .rule107(rule107[79:72]),
               .rule108(rule108[79:72]),
               .rule109(rule109[79:72]),
               .rule110(rule110[79:72]),
               .rule111(rule111[79:72]),
               .rule112(rule112[79:72]),
               .rule113(rule113[79:72]),
               .rule114(rule114[79:72]),
               .rule115(rule115[79:72]),
               .rule116(rule116[79:72]),
               .rule117(rule117[79:72]),
               .rule118(rule118[79:72]),
               .rule119(rule119[79:72]),
		.match(data9));
Row_of_RAM iRow_of_RAM10(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[87:80]),.key(key[87:80]),
		.rule0(rule0[87:80]),
		.rule1(rule1[87:80]),
		.rule2(rule2[87:80]),
		.rule3(rule3[87:80]),
		.rule4(rule4[87:80]),
		.rule5(rule5[87:80]),
		.rule6(rule6[87:80]),
		.rule7(rule7[87:80]),
		.rule8(rule8[87:80]),
		.rule9(rule9[87:80]),
		.rule10(rule10[87:80]),
		.rule11(rule11[87:80]),
		.rule12(rule12[87:80]),
		.rule13(rule13[87:80]),
		.rule14(rule14[87:80]),
                .rule15(rule15[87:80]),
                .rule16(rule16[87:80]),
                .rule17(rule17[87:80]),
                .rule18(rule18[87:80]),
                .rule19(rule19[87:80]),
                .rule20(rule20[87:80]),
                .rule21(rule21[87:80]),
                .rule22(rule22[87:80]),
                .rule23(rule23[87:80]),
                .rule24(rule24[87:80]),
                .rule25(rule25[87:80]),
                .rule26(rule26[87:80]),
                .rule27(rule27[87:80]),
                .rule28(rule28[87:80]),
                .rule29(rule29[87:80]),
                .rule30(rule30[87:80]),
                .rule31(rule31[87:80]),
                .rule32(rule32[87:80]),
                .rule33(rule33[87:80]),
               	.rule34(rule34[87:80]),
               	.rule35(rule35[87:80]),
                .rule36(rule36[87:80]),
               .rule37(rule37[87:80]),
               .rule38(rule38[87:80]),
               .rule39(rule39[87:80]),
               .rule40(rule40[87:80]),
               .rule41(rule41[87:80]),
               .rule42(rule42[87:80]),
               .rule43(rule43[87:80]),
               .rule44(rule44[87:80]),
               .rule45(rule45[87:80]),
               .rule46(rule46[87:80]),
               .rule47(rule47[87:80]),
               .rule48(rule48[87:80]),
               .rule49(rule49[87:80]),
               .rule50(rule50[87:80]),
               .rule51(rule51[87:80]),
               .rule52(rule52[87:80]),
               .rule53(rule53[87:80]),
               .rule54(rule54[87:80]),
               .rule55(rule55[87:80]),
               .rule56(rule56[87:80]),
               .rule57(rule57[87:80]),
               .rule58(rule58[87:80]),
               .rule59(rule59[87:80]),
               .rule60(rule60[87:80]),
               .rule61(rule61[87:80]),
               .rule62(rule62[87:80]),
               .rule63(rule63[87:80]),
               .rule64(rule64[87:80]),
               .rule65(rule65[87:80]),
               .rule66(rule66[87:80]),
               .rule67(rule67[87:80]),
               .rule68(rule68[87:80]),
               .rule69(rule69[87:80]),
               .rule70(rule70[87:80]),
               .rule71(rule71[87:80]),
               .rule72(rule72[87:80]),
               .rule73(rule73[87:80]),
               .rule74(rule74[87:80]),
               .rule75(rule75[87:80]),
               .rule76(rule76[87:80]),
               .rule77(rule77[87:80]),
               .rule78(rule78[87:80]),
               .rule79(rule79[87:80]),
               .rule80(rule80[87:80]),
               .rule81(rule81[87:80]),
               .rule82(rule82[87:80]),
               .rule83(rule83[87:80]),
               .rule84(rule84[87:80]),
               .rule85(rule85[87:80]),
               .rule86(rule86[87:80]),
               .rule87(rule87[87:80]),
               .rule88(rule88[87:80]),
               .rule89(rule89[87:80]),
               .rule90(rule90[87:80]),
               .rule91(rule91[87:80]),
               .rule92(rule92[87:80]),
               .rule93(rule93[87:80]),
               .rule94(rule94[87:80]),
               .rule95(rule95[87:80]),
               .rule96(rule96[87:80]),
               .rule97(rule97[87:80]),
               .rule98(rule98[87:80]),
               .rule99(rule99[87:80]),
               .rule100(rule100[87:80]),
               .rule101(rule101[87:80]),
               .rule102(rule102[87:80]),
               .rule103(rule103[87:80]),
               .rule104(rule104[87:80]),
               .rule105(rule105[87:80]),
               .rule106(rule106[87:80]),
               .rule107(rule107[87:80]),
               .rule108(rule108[87:80]),
               .rule109(rule109[87:80]),
               .rule110(rule110[87:80]),
               .rule111(rule111[87:80]),
               .rule112(rule112[87:80]),
               .rule113(rule113[87:80]),
               .rule114(rule114[87:80]),
               .rule115(rule115[87:80]),
               .rule116(rule116[87:80]),
               .rule117(rule117[87:80]),
               .rule118(rule118[87:80]),
               .rule119(rule119[87:80]),
		.match(data10));
Row_of_RAM iRow_of_RAM11(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[95:88]),.key(key[95:88]),
		.rule0(rule0[95:88]),
		.rule1(rule1[95:88]),
		.rule2(rule2[95:88]),
		.rule3(rule3[95:88]),
		.rule4(rule4[95:88]),
		.rule5(rule5[95:88]),
		.rule6(rule6[95:88]),
		.rule7(rule7[95:88]),
		.rule8(rule8[95:88]),
		.rule9(rule9[95:88]),
		.rule10(rule10[95:88]),
		.rule11(rule11[95:88]),
		.rule12(rule12[95:88]),
		.rule13(rule13[95:88]),
		.rule14(rule14[95:88]),
                .rule15(rule15[95:88]),
                .rule16(rule16[95:88]),
                .rule17(rule17[95:88]),
                .rule18(rule18[95:88]),
                .rule19(rule19[95:88]),
                .rule20(rule20[95:88]),
                .rule21(rule21[95:88]),
                .rule22(rule22[95:88]),
                .rule23(rule23[95:88]),
                .rule24(rule24[95:88]),
                .rule25(rule25[95:88]),
                .rule26(rule26[95:88]),
                .rule27(rule27[95:88]),
                .rule28(rule28[95:88]),
                .rule29(rule29[95:88]),
                .rule30(rule30[95:88]),
                .rule31(rule31[95:88]),
                .rule32(rule32[95:88]),
                .rule33(rule33[95:88]),
               	.rule34(rule34[95:88]),
               	.rule35(rule35[95:88]),
                .rule36(rule36[95:88]),
               .rule37(rule37[95:88]),
               .rule38(rule38[95:88]),
               .rule39(rule39[95:88]),
               .rule40(rule40[95:88]),
               .rule41(rule41[95:88]),
               .rule42(rule42[95:88]),
               .rule43(rule43[95:88]),
               .rule44(rule44[95:88]),
               .rule45(rule45[95:88]),
               .rule46(rule46[95:88]),
               .rule47(rule47[95:88]),
               .rule48(rule48[95:88]),
               .rule49(rule49[95:88]),
               .rule50(rule50[95:88]),
               .rule51(rule51[95:88]),
               .rule52(rule52[95:88]),
               .rule53(rule53[95:88]),
               .rule54(rule54[95:88]),
               .rule55(rule55[95:88]),
               .rule56(rule56[95:88]),
               .rule57(rule57[95:88]),
               .rule58(rule58[95:88]),
               .rule59(rule59[95:88]),
               .rule60(rule60[95:88]),
               .rule61(rule61[95:88]),
               .rule62(rule62[95:88]),
               .rule63(rule63[95:88]),
               .rule64(rule64[95:88]),
               .rule65(rule65[95:88]),
               .rule66(rule66[95:88]),
               .rule67(rule67[95:88]),
               .rule68(rule68[95:88]),
               .rule69(rule69[95:88]),
               .rule70(rule70[95:88]),
               .rule71(rule71[95:88]),
               .rule72(rule72[95:88]),
               .rule73(rule73[95:88]),
               .rule74(rule74[95:88]),
               .rule75(rule75[95:88]),
               .rule76(rule76[95:88]),
               .rule77(rule77[95:88]),
               .rule78(rule78[95:88]),
               .rule79(rule79[95:88]),
               .rule80(rule80[95:88]),
               .rule81(rule81[95:88]),
               .rule82(rule82[95:88]),
               .rule83(rule83[95:88]),
               .rule84(rule84[95:88]),
               .rule85(rule85[95:88]),
               .rule86(rule86[95:88]),
               .rule87(rule87[95:88]),
               .rule88(rule88[95:88]),
               .rule89(rule89[95:88]),
               .rule90(rule90[95:88]),
               .rule91(rule91[95:88]),
               .rule92(rule92[95:88]),
               .rule93(rule93[95:88]),
               .rule94(rule94[95:88]),
               .rule95(rule95[95:88]),
               .rule96(rule96[95:88]),
               .rule97(rule97[95:88]),
               .rule98(rule98[95:88]),
               .rule99(rule99[95:88]),
               .rule100(rule100[95:88]),
               .rule101(rule101[95:88]),
               .rule102(rule102[95:88]),
               .rule103(rule103[95:88]),
               .rule104(rule104[95:88]),
               .rule105(rule105[95:88]),
               .rule106(rule106[95:88]),
               .rule107(rule107[95:88]),
               .rule108(rule108[95:88]),
               .rule109(rule109[95:88]),
               .rule110(rule110[95:88]),
               .rule111(rule111[95:88]),
               .rule112(rule112[95:88]),
               .rule113(rule113[95:88]),
               .rule114(rule114[95:88]),
               .rule115(rule115[95:88]),
               .rule116(rule116[95:88]),
               .rule117(rule117[95:88]),
               .rule118(rule118[95:88]),
               .rule119(rule119[95:88]),
		.match(data11));
Row_of_RAM iRow_of_RAM13(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[103:96]),.key(key[103:96]),
		.rule0(rule0[103:96]),
		.rule1(rule1[103:96]),
		.rule2(rule2[103:96]),
		.rule3(rule3[103:96]),
		.rule4(rule4[103:96]),
		.rule5(rule5[103:96]),
		.rule6(rule6[103:96]),
		.rule7(rule7[103:96]),
		.rule8(rule8[103:96]),
		.rule9(rule9[103:96]),
		.rule10(rule10[103:96]),
		.rule11(rule11[103:96]),
		.rule12(rule12[103:96]),
		.rule13(rule13[103:96]),
		.rule14(rule14[103:96]),
                .rule15(rule15[103:96]),
                .rule16(rule16[103:96]),
                .rule17(rule17[103:96]),
                .rule18(rule18[103:96]),
                .rule19(rule19[103:96]),
                .rule20(rule20[103:96]),
                .rule21(rule21[103:96]),
                .rule22(rule22[103:96]),
                .rule23(rule23[103:96]),
                .rule24(rule24[103:96]),
                .rule25(rule25[103:96]),
                .rule26(rule26[103:96]),
                .rule27(rule27[103:96]),
                .rule28(rule28[103:96]),
                .rule29(rule29[103:96]),
                .rule30(rule30[103:96]),
                .rule31(rule31[103:96]),
                .rule32(rule32[103:96]),
                .rule33(rule33[103:96]),
               	.rule34(rule34[103:96]),
               	.rule35(rule35[103:96]),
                .rule36(rule36[103:96]),
               .rule37(rule37[103:96]),
               .rule38(rule38[103:96]),
               .rule39(rule39[103:96]),
               .rule40(rule40[103:96]),
               .rule41(rule41[103:96]),
               .rule42(rule42[103:96]),
               .rule43(rule43[103:96]),
               .rule44(rule44[103:96]),
               .rule45(rule45[103:96]),
               .rule46(rule46[103:96]),
               .rule47(rule47[103:96]),
               .rule48(rule48[103:96]),
               .rule49(rule49[103:96]),
               .rule50(rule50[103:96]),
               .rule51(rule51[103:96]),
               .rule52(rule52[103:96]),
               .rule53(rule53[103:96]),
               .rule54(rule54[103:96]),
               .rule55(rule55[103:96]),
               .rule56(rule56[103:96]),
               .rule57(rule57[103:96]),
               .rule58(rule58[103:96]),
               .rule59(rule59[103:96]),
               .rule60(rule60[103:96]),
               .rule61(rule61[103:96]),
               .rule62(rule62[103:96]),
               .rule63(rule63[103:96]),
               .rule64(rule64[103:96]),
               .rule65(rule65[103:96]),
               .rule66(rule66[103:96]),
               .rule67(rule67[103:96]),
               .rule68(rule68[103:96]),
               .rule69(rule69[103:96]),
               .rule70(rule70[103:96]),
               .rule71(rule71[103:96]),
               .rule72(rule72[103:96]),
               .rule73(rule73[103:96]),
               .rule74(rule74[103:96]),
               .rule75(rule75[103:96]),
               .rule76(rule76[103:96]),
               .rule77(rule77[103:96]),
               .rule78(rule78[103:96]),
               .rule79(rule79[103:96]),
               .rule80(rule80[103:96]),
               .rule81(rule81[103:96]),
               .rule82(rule82[103:96]),
               .rule83(rule83[103:96]),
               .rule84(rule84[103:96]),
               .rule85(rule85[103:96]),
               .rule86(rule86[103:96]),
               .rule87(rule87[103:96]),
               .rule88(rule88[103:96]),
               .rule89(rule89[103:96]),
               .rule90(rule90[103:96]),
               .rule91(rule91[103:96]),
               .rule92(rule92[103:96]),
               .rule93(rule93[103:96]),
               .rule94(rule94[103:96]),
               .rule95(rule95[103:96]),
               .rule96(rule96[103:96]),
               .rule97(rule97[103:96]),
               .rule98(rule98[103:96]),
               .rule99(rule99[103:96]),
               .rule100(rule100[103:96]),
               .rule101(rule101[103:96]),
               .rule102(rule102[103:96]),
               .rule103(rule103[103:96]),
               .rule104(rule104[103:96]),
               .rule105(rule105[103:96]),
               .rule106(rule106[103:96]),
               .rule107(rule107[103:96]),
               .rule108(rule108[103:96]),
               .rule109(rule109[103:96]),
               .rule110(rule110[103:96]),
               .rule111(rule111[103:96]),
               .rule112(rule112[103:96]),
               .rule113(rule113[103:96]),
               .rule114(rule114[103:96]),
               .rule115(rule115[103:96]),
               .rule116(rule116[103:96]),
               .rule117(rule117[103:96]),
               .rule118(rule118[103:96]),
               .rule119(rule119[103:96]),
		.match(data12));

assign i_data = data0 & data1 & data2 & data3 & data4 & data5 & data6 & data7 & data8 & data9 & data10 & data11 & data12;

always @(i_data)  begin
	if(~resetn) begin
          result <= 120'b0;
	end else
         result <= i_data;
   
end



endmodule





