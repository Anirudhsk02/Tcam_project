module Row_of_RAM(input write_clk,
                input wren,
                input readen,
                input [7:0] wr_addr,
                input [7:0] key, // key = read_addr
                input [7:0] rule0,
                input [7:0] rule1,
                input [7:0] rule2,
                input [7:0] rule3,
                input [7:0] rule4,
                input [7:0] rule5,
                input [7:0] rule6,
                input [7:0] rule7,
                input [7:0] rule8,
                input [7:0] rule9,
                input [7:0] rule10,
                input [7:0] rule11,
                input [7:0] rule12,
                input [7:0] rule13,
                input [7:0] rule14,
                input [7:0] rule15,
                input [7:0] rule16,
                input [7:0] rule17,
                input [7:0] rule18,
                input [7:0] rule19,
                input [7:0] rule20,
                input [7:0] rule21,
                input [7:0] rule22,
                input [7:0] rule23,
                input [7:0] rule24,
                input [7:0] rule25,
                input [7:0] rule26,
                input [7:0] rule27,
                input [7:0] rule28,
                input [7:0] rule29,
                input [7:0] rule30,
                input [7:0] rule31,
                input [7:0] rule32,
                input [7:0] rule33,
               input [7:0] rule34,
               input [7:0] rule35,
               input [7:0] rule36,
               input [7:0] rule37,
               input [7:0] rule38,
               input [7:0] rule39,
               input [7:0] rule40,
               input [7:0] rule41,
               input [7:0] rule42,
               input [7:0] rule43,
               input [7:0] rule44,
               input [7:0] rule45,
               input [7:0] rule46,
               input [7:0] rule47,
               input [7:0] rule48,
               input [7:0] rule49,
               input [7:0] rule50,
               input [7:0] rule51,
               input [7:0] rule52,
               input [7:0] rule53,
               input [7:0] rule54,
               input [7:0] rule55,
               input [7:0] rule56,
               input [7:0] rule57,
               input [7:0] rule58,
               input [7:0] rule59,
               input [7:0] rule60,
               input [7:0] rule61,
               input [7:0] rule62,
               input [7:0] rule63,
               input [7:0] rule64,
               input [7:0] rule65,
               input [7:0] rule66,
               input [7:0] rule67,
               input [7:0] rule68,
               input [7:0] rule69,
               input [7:0] rule70,
               input [7:0] rule71,
               input [7:0] rule72,
               input [7:0] rule73,
               input [7:0] rule74,
               input [7:0] rule75,
               input [7:0] rule76,
               input [7:0] rule77,
               input [7:0] rule78,
               input [7:0] rule79,
               input [7:0] rule80,
               input [7:0] rule81,
               input [7:0] rule82,
               input [7:0] rule83,
               input [7:0] rule84,
               input [7:0] rule85,
               input [7:0] rule86,
               input [7:0] rule87,
               input [7:0] rule88,
               input [7:0] rule89,
               input [7:0] rule90,
               input [7:0] rule91,
               input [7:0] rule92,
               input [7:0] rule93,
               input [7:0] rule94,
               input [7:0] rule95,
               input [7:0] rule96,
               input [7:0] rule97,
               input [7:0] rule98,
               input [7:0] rule99,
               input [7:0] rule100,
               input [7:0] rule101,
               input [7:0] rule102,
               input [7:0] rule103,
               input [7:0] rule104,
               input [7:0] rule105,
               input [7:0] rule106,
               input [7:0] rule107,
               input [7:0] rule108,
               input [7:0] rule109,
               input [7:0] rule110,
               input [7:0] rule111,
               input [7:0] rule112,
               input [7:0] rule113,
               input [7:0] rule114,
               input [7:0] rule115,
               input [7:0] rule116,
                input [7:0] rule117,
                input [7:0] rule118,
                input [7:0] rule119,
                

                output  [119:0] match
        );


             RAM_8bit iRAM_8bit1(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule0[7:0]),.rule1(rule1[7:0]),.rule2(rule2[7:0]),.rule3(rule3[7:0]),.rule4(rule4[7:0]),.rule5(rule5[7:0]),.rule6(rule6[7:0]),.rule7(rule7[7:0]),.match(match[7:0]));
             RAM_8bit iRAM_8bit2(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule8[7:0]),.rule1(rule9[7:0]),.rule2(rule10[7:0]),.rule3(rule11[7:0]),.rule4(rule12[7:0]),.rule5(rule13[7:0]),.rule6(rule14[7:0]),.rule7(rule15[7:0]),.match(match[15:8]));
             RAM_8bit iRAM_8bit3(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule16[7:0]),.rule1(rule17[7:0]),.rule2(rule18[7:0]),.rule3(rule19[7:0]),.rule4(rule20[7:0]),.rule5(rule21[7:0]),.rule6(rule22[7:0]),.rule7(rule23[7:0]),.match(match[23:16]));
             RAM_8bit iRAM_8bit4(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule24[7:0]),.rule1(rule25[7:0]),.rule2(rule26[7:0]),.rule3(rule27[7:0]),.rule4(rule28[7:0]),.rule5(rule29[7:0]),.rule6(rule30[7:0]),.rule7(rule31[7:0]),.match(match[31:24]));
             RAM_8bit iRAM_8bit5(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule32[7:0]),.rule1(rule33[7:0]),.rule2(rule34[7:0]),.rule3(rule35[7:0]),.rule4(rule36[7:0]),.rule5(rule37[7:0]),.rule6(rule38[7:0]),.rule7(rule39[7:0]),.match(match[39:32]));
             RAM_8bit iRAM_8bit6(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule40[7:0]),.rule1(rule41[7:0]),.rule2(rule42[7:0]),.rule3(rule43[7:0]),.rule4(rule44[7:0]),.rule5(rule45[7:0]),.rule6(rule46[7:0]),.rule7(rule47[7:0]),.match(match[47:40]));
             RAM_8bit iRAM_8bit7(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule48[7:0]),.rule1(rule49[7:0]),.rule2(rule50[7:0]),.rule3(rule51[7:0]),.rule4(rule52[7:0]),.rule5(rule53[7:0]),.rule6(rule54[7:0]),.rule7(rule55[7:0]),.match(match[55:48]));
             RAM_8bit iRAM_8bit8(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule56[7:0]),.rule1(rule57[7:0]),.rule2(rule58[7:0]),.rule3(rule59[7:0]),.rule4(rule60[7:0]),.rule5(rule61[7:0]),.rule6(rule62[7:0]),.rule7(rule63[7:0]),.match(match[63:56]));
             RAM_8bit iRAM_8bit9(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule64[7:0]),.rule1(rule65[7:0]),.rule2(rule66[7:0]),.rule3(rule67[7:0]),.rule4(rule68[7:0]),.rule5(rule69[7:0]),.rule6(rule70[7:0]),.rule7(rule71[7:0]),.match(match[71:64]));
             RAM_8bit iRAM_8bit10(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule72[7:0]),.rule1(rule73[7:0]),.rule2(rule74[7:0]),.rule3(rule75[7:0]),.rule4(rule76[7:0]),.rule5(rule77[7:0]),.rule6(rule78[7:0]),.rule7(rule79[7:0]),.match(match[79:72]));
             RAM_8bit iRAM_8bit11(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule80[7:0]),.rule1(rule81[7:0]),.rule2(rule82[7:0]),.rule3(rule83[7:0]),.rule4(rule84[7:0]),.rule5(rule85[7:0]),.rule6(rule86[7:0]),.rule7(rule87[7:0]),.match(match[87:80]));
             RAM_8bit iRAM_8bit12(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule88[7:0]),.rule1(rule89[7:0]),.rule2(rule90[7:0]),.rule3(rule91[7:0]),.rule4(rule92[7:0]),.rule5(rule93[7:0]),.rule6(rule94[7:0]),.rule7(rule95[7:0]),.match(match[95:88]));
             RAM_8bit iRAM_8bit13(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule96[7:0]),.rule1(rule97[7:0]),.rule2(rule98[7:0]),.rule3(rule99[7:0]),.rule4(rule100[7:0]),.rule5(rule101[7:0]),.rule6(rule102[7:0]),.rule7(rule103[7:0]),.match(match[103:96]));
             RAM_8bit iRAM_8bit14(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule104[7:0]),.rule1(rule105[7:0]),.rule2(rule106[7:0]),.rule3(rule107[7:0]),.rule4(rule108[7:0]),.rule5(rule109[7:0]),.rule6(rule110[7:0]),.rule7(rule111[7:0]),.match(match[111:104]));
             RAM_8bit iRAM_8bit15(.write_clk(write_clk),.wren(wren),.readen(readen),.wr_addr(wr_addr[7:0]),.key(key[7:0]),.rule0(rule112[7:0]),.rule1(rule113[7:0]),.rule2(rule114[7:0]),.rule3(rule115[7:0]),.rule4(rule116[7:0]),.rule5(rule117[7:0]),.rule6(rule118[7:0]),.rule7(rule119[7:0]),.match(match[119:112]));



        endmodule
